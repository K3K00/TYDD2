library verilog;
use verilog.vl_types.all;
entity restador_completo_vlg_check_tst is
    port(
        o_bout          : in     vl_logic;
        o_rout          : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end restador_completo_vlg_check_tst;
